.title KiCad schematic
.include "models/C2012C0G1H153J085AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C3216X7R1H105K160AB_p.mod"
.include "models/MJD31C.spice.txt"
.include "models/XPE_SPICE.lib"
.include "models/max16823.lib"
XU3 /DIMM /DIMM /DIMM /LEDGOOD VCC /LGC /REG 0 /SENSE3 /SENSE2 /SENSE1 /CHN3 /CHN2 /CHN1 MAX16823
XU2 VCC 0 C2012X7R2A104K125AA_p
R2 /SENSE1 0 {Rsense}
R3 /SENSE2 0 {Rsense}
R4 /SENSE3 0 {Rsense}
R1 /REG /LEDGOOD 10k
XU1 /REG 0 C2012X7R2A104K125AA_p
V1 VCC 0 {Vin}
V2 /DIMM 0 PULSE(0 {vpul} 0 {tr} {tf} {duty} {cycle})
XU4 /LGC 0 C2012C0G1H153J085AA_p
Q1 VCC /CHN1 /G_1 MJD31C
R5 /CHN1 0 {Rpd}
R6 /CHN2 0 {Rpd}
R7 /CHN3 0 {Rpd}
D9 /R_3 /SENSE3 XLampXPEred
D8 /B_3 /SENSE2 XLampXPEblue
D7 /G_3 /SENSE1 XLampXPEgreen
D5 /R_1 /R_2 XLampXPEred
D3 /B_1 /B_2 XLampXPEblue
D6 /R_2 /R_3 XLampXPEred
D4 /B_2 /B_3 XLampXPEblue
D2 /G_2 /G_3 XLampXPEgreen
D1 /G_1 /G_2 XLampXPEgreen
XU5 0 /G_1 C3216X7R1H105K160AB_p
XU6 0 /B_1 C3216X7R1H105K160AB_p
XU7 0 /R_1 C3216X7R1H105K160AB_p
XU8 0 VCC C3216X7R1H105K160AB_p
Q2 VCC /CHN2 /B_1 MJD31C
Q3 VCC /CHN3 /R_1 MJD31C
.end
